// 32_bit_unsigned_adder